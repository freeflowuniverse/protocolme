module system

pub struct Tag {
pub mut:
	name        string
	value		string 
}

