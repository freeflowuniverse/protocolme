module objtypes


fn test_1() {

	mut o:=get(1,"") or {panic(err)}
	println(o)

	println(o.json())
	
	panic("s")

}