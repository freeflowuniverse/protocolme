module people

[heap]
pub struct Country { 
pub mut:
	name  		string
	code2 		string
	code3 		string
	nr    		int
	vat_percent int = 20 //0-100
}


