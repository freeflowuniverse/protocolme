module system


[heap]
struct Remark {
pub mut:
	content string
	time    OurTime
	author  string //smartid to twin.person 
}

