module backoffice

//import freeflowuniverse.backoffice.organization
//import freeflowuniverse.crystallib.texttools

// TODO circle_add

// TODO circle_end
/*
// Find a specific Circle
pub fn (mut data Data) circle_find(circle_name string) ?&organization.Circle {
	shortname := texttools.name_fix_no_underscore_no_ext(circle_name)

	if shortname in data.circles {
		return data.circles[shortname]
	}
	return error('Could not find circle with name: $shortname')
}
*/