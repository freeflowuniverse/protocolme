module planner

[heap]
pub struct Tags {
pub mut:
	tags []Tag
}

pub struct Tag {
pub mut:
	name        string
	value		string 
}

